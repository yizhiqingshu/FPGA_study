library verilog;
use verilog.vl_types.all;
entity block_nblock_db is
end block_nblock_db;
