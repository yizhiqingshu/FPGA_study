library verilog;
use verilog.vl_types.all;
entity BCD_Counter_top_tb is
end BCD_Counter_top_tb;
